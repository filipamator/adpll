fp_int32_inst : fp_int32 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
