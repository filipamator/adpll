fp_mult_inst : fp_mult PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
